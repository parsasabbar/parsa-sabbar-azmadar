module pcadder(input[63:0]a,output[63:0] b);
  fa64b p0(64'h0000000000000004,a,1'b0,b,);
endmodule


